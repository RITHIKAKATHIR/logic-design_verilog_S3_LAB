module xor_gatelevel(y,a,b);
output y;
input a,b;
xor(y,a,b);

endmodule 