module dflipflop_assn(d, clk, enable, reset, out);
input d, clk, enable, reset;
output out;
reg out;
always @ (posedge clk or posedge reset) begin
    if (reset)
      out = 0;
    else
      if (enable)
        out = d;
 end
endmodule
