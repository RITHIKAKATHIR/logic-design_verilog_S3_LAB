module xnor_gatelevel(y,a,b);
 
input a,b;
output y;

xnor(y,a,b);

endmodule 