module nand_gatelevel(y,a,b);

input a,b;
output y;

nand(y,a,b);

endmodule

