module nor_gatelevel(y,a,b);
input a,b;
output y;

nor(y,a,b);
endmodule 
