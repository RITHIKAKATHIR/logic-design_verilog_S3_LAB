module test_1tb;

reg a,b,c;
wire y;

test_1 obj(a,b,c,y);

initial 
 begin 
    a=0;b=0;c=0;
#10 a=0;b=0;c=1;
#10 a=0;b=1;c=0;
#10 a=0;b=1;c=1;
#10 a=1;b=0;c=0;
#10 a=1;b=0;c=1;
#10 a=1;b=1;c=0;
#10 a=1;b=1;c=1;
 end
 


endmodule
