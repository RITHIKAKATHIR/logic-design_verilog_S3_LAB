module nand_input_gatelevel(out,a,b,c,d,e,f,g,h);
input a,b,c,d,e,f,g,h;
output out;
nand(out,a,b,c,d,e,f,g,h);
endmodule 
