module nor_input_gatelevel(y,a,b,c,d,e,f,g,h);
input a,b,c,d,e,f,g,h;
output y;
nor(y,a,b,c,d,e,f,g,h);

endmodule
