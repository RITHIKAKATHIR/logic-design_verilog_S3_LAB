module carrysel32_tb;
reg[31:0] sum;
reg carryout;
wire in1[0],in2[0] , in1[1],in2[1] , in1[2],in2[2] , in1[3],in2[3] , in1[4],in2[4] ,in1[5],in2[5] , in1[6],in2[6] , in1[7],in2[7]  ,in1[8],in2[8] , in1[9],in2[9] , in1[10],in2[10] , in1[11],in2[11] , in1[12],in2[12] , in1[13],in2[13] , in1[14],in2[14] , in1[15],in2[15] , in1[16],in2[16] , in1[17],in2[17] , in1[18],in2[18] , in1[19],in2[19]  ,in1[20],in2[20] , in1[21],in2[21]  ,in1[22],in2[22],  in1[23],in2[23]  ,in1[24],in2[24],  in1[25],in2[25],  in1[26],in2[26] , in1[27],in2[27] , in1[28],in2[28] ,in1[29],in2[29], in1[30],in2[30],in1[31],in2[31] ;
carryselectadder32_datafow obj(.sum(sum),.in1(in1),.in2(in2),.carryout(carryout));
initial 
  begin 
    assign in1[0]=0; in1[1]=0; in1[2]=0; in1[3]=0; in1[4]=0; in1[5]=0; in1[6]=0; in1[7]=0; in1[8]=0; in1[9]=0; in1[10]=0; in1[11]=0; in1[12]=0; in1[13]=0; in1[14]=0; in1[15]=0; in1[16]=0; in1[17]=0; in1[18]=0; in1[19]=0; in1[20]=0; in1[21]=0; in1[22]=0; in1[23]=0; in1[24]=0; in1[25]=0; in1[26]=0; in1[27]=0; in1[28]=0; in1[29]=0; in1[30]=0; in1[31]=0; 
   assign   in2[0]=0; in2[1]=0; in2[2]=0; in2[3]=0; in2[4]=0; in2[5]=0; in2[6]=0; in2[7]=0; in2[8]=0; in2[9]=0; in2[10]=0; in2[11]=0; in2[12]=0; in2[13]=0; in2[14]=0; in2[15]=0; in2[16]=0; in2[17]=0; in2[18]=0; in2[19]=0; in2[20]=0; in2[21]=0; in2[22]=0; in2[23]=0; in2[24]=0; in2[25]=0; in2[26]=0; in2[27]=0; in2[28]=0; in2[29]=0; in2[30]=0; in2[31]=0; 


   #10
assign	in1[0]=1; in1[1]=1; in1[2]=1; in1[3]=1; in1[4]=1; in1[5]=1; in1[6]=1; in1[7]=1; in1[8]=1; in1[9]=1; in1[10]=1; in1[11]=1; in1[12]=1; in1[13]=1; in1[14]=1; in1[15]=1; in1[16]=1; in1[17]=1; in1[18]=1; in1[19]=1; in1[20]=1; in1[21]=1; in1[22]=1; in1[23]=1; in1[24]=1; in1[25]=1; in1[26]=1; in1[27]=1; in1[28]=1; in1[29]=1; in1[30]=1; in1[31]=1; 
 assign   in2[0]=0; in2[1]=0; in2[2]=0; in2[3]=0; in2[4]=0; in2[5]=0; in2[6]=0; in2[7]=0; in2[8]=0; in2[9]=0; in2[10]=0; in2[11]=0; in2[12]=0; in2[13]=0; in2[14]=0; in2[15]=0; in2[16]=0; in2[17]=0; in2[18]=0; in2[19]=0; in2[20]=0; in2[21]=0; in2[22]=0; in2[23]=0; in2[24]=0; in2[25]=0; in2[26]=0; in2[27]=0; in2[28]=0; in2[29]=0; in2[30]=0; in2[31]=0; 

   #10
assign	in1[0]=0; in1[1]=0; in1[2]=0; in1[3]=0; in1[4]=0; in1[5]=0; in1[6]=0; in1[7]=0; in1[8]=0; in1[9]=0; in1[10]=0; in1[11]=0; in1[12]=0; in1[13]=0; in1[14]=0; in1[15]=0; in1[16]=0; in1[17]=0; in1[18]=0; in1[19]=0; in1[20]=0; in1[21]=0; in1[22]=0; in1[23]=0; in1[24]=0; in1[25]=0; in1[26]=0; in1[27]=0; in1[28]=0; in1[29]=0; in1[30]=0; in1[31]=0; 

assign	in2[0]=1; in2[1]=1; in2[2]=1; in2[3]=1; in2[4]=1; in2[5]=1; in2[6]=1; in2[7]=1; in2[8]=1; in2[9]=1; in2[10]=1; in2[11]=1; in2[12]=1; in2[13]=1; in2[14]=1; in2[15]=1; in2[16]=1; in2[17]=1; in2[18]=1; in2[19]=1; in2[20]=1; in2[21]=1; in2[22]=1; in2[23]=1; in2[24]=1; in2[25]=1; in2[26]=1; in2[27]=1; in2[28]=1; in2[29]=1; in2[30]=1; in2[31]=1; 
   #10
assign	in1[0]=1; in1[1]=1; in1[2]=1; in1[3]=1; in1[4]=1; in1[5]=1; in1[6]=1; in1[7]=1; in1[8]=1; in1[9]=1; in1[10]=1; in1[11]=1; in1[12]=1; in1[13]=1; in1[14]=1; in1[15]=1; in1[16]=1; in1[17]=1; in1[18]=1; in1[19]=1; in1[20]=1; in1[21]=1; in1[22]=1; in1[23]=1; in1[24]=1; in1[25]=1; in1[26]=1; in1[27]=1; in1[28]=1; in1[29]=1; in1[30]=1; in1[31]=1; 
assign   in2[0]=1; in2[1]=1; in2[2]=1; in2[3]=1; in2[4]=1; in2[5]=1; in2[6]=1; in2[7]=1; in2[8]=1; in2[9]=1; in2[10]=1; in2[11]=1; in2[12]=1; in2[13]=1; in2[14]=1; in2[15]=1; in2[16]=1; in2[17]=1; in2[18]=1; in2[19]=1; in2[20]=1; in2[21]=1; in2[22]=1; in2[23]=1; in2[24]=1; in2[25]=1; in2[26]=1; in2[27]=1; in2[28]=1; in2[29]=1; in2[30]=1; in2[31]=1; 

  
 end
  
endmodule
