module add_gate_gatelevel(y,a,b);

input a;
input b;
output y;

and(y,a,b);
endmodule 