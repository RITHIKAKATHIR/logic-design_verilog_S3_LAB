module inverter_gate_level(out,in);
output out;
input in;
not(out,in);

endmodule 