module or_gate_gatelevel(y,a,b);
input a,b;
output y;

or(y,a,b);

endmodule
