module carry_select_adder()